module Pratica01 (
	output 	[7:0] LED
);

assign LED = 'h55;

endmodule
